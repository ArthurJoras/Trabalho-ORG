----------------------------------------------------------------------------------
-- Company: UERGS
-- Engineer: Arthur Joras && Artur de Camargo .
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.ALL;

entity memory is
	port(		
        clk                 : in  std_logic;
        escrita             : in  std_logic;
		leitura             : in  std_logic;
        rst_n               : in  std_logic;        
        entrada_memoria     : in  std_logic_vector(15 downto 0);
        endereco_memoria    : in  std_logic_vector(7  downto 0);
        saida_memoria       : out std_logic_vector(15 downto 0)
	);
        
end memory;

architecture rtl of memory is

	-- 256 words of 2 bytes (16 bits)
	subtype palavra is std_logic_vector(15 downto 0);
	type memory is array (0 to 255) of palavra;
	signal mem : memory;
	
begin 

process(clk)	
begin
			
	if(rst_n = '1') then
		--  reset memory when rst_n = 1  
		mem(0)    <= "0000000000000000"; 
		mem(1)    <= "0000000000000000";
		mem(2)    <= "0000000000000000";
		mem(3)    <= "0000000000000000";
		mem(4)    <= "0000000000000000";
		mem(5)    <= "0000000000000000"; 
		mem(6)    <= "0000000000000000";
		mem(7)    <= "0000000000000000";
		mem(8)    <= "0000000000000000";
		mem(9)    <= "0000000000000000";
		mem(10)   <= "0000000000000000";
		mem(11)   <= "0000000000000000";
		mem(12)   <= "0000000000000000";
		mem(13)   <= "0000000000000000";
		mem(14)   <= "0000000000000000";
		mem(15)   <= "0000000000000000"; 
		mem(16)   <= "0000000000000000"; 
		mem(17)   <= "0000000000000000"; 
		mem(18)   <= "0000000000000000"; 
		mem(19)   <= "0000000000000000"; 
		mem(20)   <= "0000000000000000";
		mem(21)   <= "0000000000000000"; 
		mem(22)   <= "0000000000000000";
		mem(23)   <= "0000000000000000";
		mem(24)   <= "0000000000000000"; 
		mem(25)   <= "0000000000000000"; 
		mem(26)   <= "0000000000000000"; 
		mem(27)   <= "0000000000000000";      
		mem(28)   <= "0000000000000000"; 
		mem(29)   <= "0000000000000000"; 
		mem(30)   <= "0000000000000000"; 
		mem(31)   <= "0000000000000000"; 
		mem(32)   <= "0000000000000000";  
		mem(33)   <= "0000000000000000"; 
		mem(34)   <= "0000000000000000"; 
		mem(35)   <= "0000000000000000";
		mem(36)   <= "0000000000000000";
		mem(37)   <= "0000000000000000";
		mem(38)   <= "0000000000000000";
		mem(39)   <= "0000000000000000";
		mem(40)   <= "0000000000000000";
		mem(41)   <= "0000000000000000";
		mem(42)   <= "0000000000000000";
		mem(43)   <= "0000000000000000";
		mem(44)   <= "0000000000000000";
		mem(45)   <= "0000000000000000";
		mem(46)   <= "0000000000000000";
		mem(47)   <= "0000000000000000";
		mem(48)   <= "0000000000000000";
		mem(49)   <= "0000000000000000";
		mem(50)   <= "0000000000000000";
		mem(51)   <= "0000000000000000"; 
		mem(52)   <= "0000000000000000";
		mem(53)   <= "0000000000000000";
		mem(54)   <= "0000000000000000";
		mem(55)   <= "0000000000000000";
		mem(56)   <= "0000000000000000";
		mem(57)   <= "0000000000000000";
		mem(58)   <= "0000000000000000";
		mem(59)   <= "0000000000000000";
		mem(60)   <= "0000000000000000";
		mem(61)   <= "0000000000000000";
		mem(62)   <= "0000000000000000";
		mem(63)   <= "0000000000000000";
		mem(64)   <= "0000000000000000";
		mem(65)   <= "0000000000000000";
		mem(66)   <= "0000000000000000"; 
		mem(67)   <= "0000000000000000";
		mem(68)   <= "0000000000000000"; 
		mem(69)   <= "0000000000000000";
		mem(70)   <= "0000000000000000";
		mem(71)   <= "0000000000000000";
		mem(72)   <= "0000000000000000";
		mem(73)   <= "0000000000000000";
		mem(74)   <= "0000000000000000"; 
		mem(75)   <= "0000000000000000";
		mem(76)   <= "0000000000000000";
		mem(77)   <= "0000000000000000";
		mem(78)   <= "0000000000000000"; 
		mem(79)   <= "0000000000000000";
		mem(80)   <= "0000000000000000"; 
		mem(81)   <= "0000000000000000";
		mem(82)   <= "0000000000000000";  
		mem(83)   <= "0000000000000000";
		mem(84)   <= "0000000000000000";
		mem(85)   <= "0000000000000000";
		mem(86)   <= "0000000000000000";
		mem(87)   <= "0000000000000000";
		mem(88)   <= "0000000000000000";
		mem(89)   <= "0000000000000000";
		mem(90)   <= "0000000000000000";
		mem(91)   <= "0000000000000000";
		mem(92)   <= "0000000000000000";
		mem(93)   <= "0000000000000000";
		mem(94)   <= "0000000000000000";
		mem(95)   <= "0000000000000000";
		mem(96)   <= "0000000000000000";
		mem(97)   <= "0000000000000000";
		mem(98)   <= "0000000000000000";
		mem(99)   <= "0000000000000000";
		mem(100)  <= "0000000000000000"; 
		mem(101)  <= "0000000000000000";
		mem(102)  <= "0000000000000000"; 
		mem(103)  <= "0000000000000000";
		mem(104)  <= "0000000000000000";
		mem(105)  <= "0000000000000000";
		mem(106)  <= "0000000000000000";
		mem(107)  <= "0000000000000000";
		mem(108)  <= "0000000000000000";
		mem(109)  <= "0000000000000000";
		mem(110)  <= "0000000000000000";
		mem(111)  <= "0000000000000000";
		mem(112)  <= "0000000000000000";
		mem(113)  <= "0000000000000000";
		mem(114)  <= "0000000000000000";
		mem(115)  <= "0000000000000000";
		mem(116)  <= "0000000000000000";
		mem(117)  <= "0000000000000000";
		mem(118)  <= "0000000000000000";
		mem(119)  <= "0000000000000000";
		mem(120)  <= "0000000000000000";
		mem(121)  <= "0000000000000000";
		mem(122)  <= "0000000000000000";
		mem(123)  <= "0000000000000000";
		mem(124)  <= "0000000000000000";
		mem(125)  <= "0000000000000000";
		mem(126)  <= "0000000000000000";
		mem(127)  <= "0000000000000000";
		mem(128)  <= "0000000000000000";
		mem(129)  <= "0000000000000000"; 
		mem(130)  <= "0000000000000000"; 
		mem(131)  <= "0000000000000000";
		mem(132)  <= "0000000000000000";
		mem(133)  <= "0000000000000000";
		mem(134)  <= "0000000000000000";
		mem(135)  <= "0000000000000000";
		mem(136)  <= "0000000000000000";
		mem(137)  <= "0000000000000000";
		mem(138)  <= "0000000000000000";
		mem(139)  <= "0000000000000000";
		mem(140)  <= "0000000000000000";
		mem(141)  <= "0000000000000000";
		mem(142)  <= "0000000000000000";
		mem(143)  <= "0000000000000000";
		mem(144)  <= "0000000000000000";
		mem(145)  <= "0000000000000000";
		mem(146)  <= "0000000000000000";
		mem(147)  <= "0000000000000000";
		mem(148)  <= "0000000000000000";
		mem(149)  <= "0000000000000000";
		mem(150)  <= "0000000000000000";
		mem(151)  <= "0000000000000000";
		mem(152)  <= "0000000000000000";
		mem(153)  <= "0000000000000000";
		mem(154)  <= "0000000000000000";
		mem(155)  <= "0000000000000000";
		mem(156)  <= "0000000000000000";
		mem(157)  <= "0000000000000000";
		mem(158)  <= "0000000000000000";
		mem(159)  <= "0000000000000000";
		mem(160)  <= "0000000000000000";
		mem(161)  <= "0000000000000000";
		mem(162)  <= "0000000000000000";
		mem(163)  <= "0000000000000000";
		mem(164)  <= "0000000000000000";
		mem(165)  <= "0000000000000000";
		mem(166)  <= "0000000000000000";
		mem(167)  <= "0000000000000000";
		mem(168)  <= "0000000000000000";
		mem(169)  <= "0000000000000000";
		mem(170)  <= "0000000000000000";
		mem(171)  <= "0000000000000000";
		mem(172)  <= "0000000000000000";
		mem(173)  <= "0000000000000000";
		mem(174)  <= "0000000000000000";
		mem(175)  <= "0000000000000000";
		mem(176)  <= "0000000000000000";
		mem(177)  <= "0000000000000000";
		mem(178)  <= "0000000000000000";
		mem(179)  <= "0000000000000000";
		mem(180)  <= "0000000000000000";
		mem(181)  <= "0000000000000000";
		mem(182)  <= "0000000000000000";
		mem(183)  <= "0000000000000000";
		mem(184)  <= "0000000000000000";
		mem(185)  <= "0000000000000000";
		mem(186)  <= "0000000000000000";
		mem(187)  <= "0000000000000000";
		mem(188)  <= "0000000000000000";
		mem(189)  <= "0000000000000000";
		mem(190)  <= "0000000000000000";
		mem(191)  <= "0000000000000000";
		mem(192)  <= "0000000000000000";
		mem(193)  <= "0000000000000000";
		mem(194)  <= "0000000000000000";
		mem(195)  <= "0000000000000000";
		mem(196)  <= "0000000000000000";
		mem(197)  <= "0000000000000000";
		mem(198)  <= "0000000000000000";
		mem(199)  <= "0000000000000000";
		mem(200)  <= "0000000000000000";
		mem(201)  <= "0000000000000000";
		mem(202)  <= "0000000000000000";
		mem(203)  <= "0000000000000000";
		mem(204)  <= "0000000000000000";
		mem(205)  <= "0000000000000000";
		mem(206)  <= "0000000000000000";
		mem(207)  <= "0000000000000000";
		mem(208)  <= "0000000000000000";
		mem(209)  <= "0000000000000000";
		mem(210)  <= "0000000000000000";
		mem(211)  <= "0000000000000000";
		mem(212)  <= "0000000000000000";
		mem(213)  <= "0000000000000000";
		mem(214)  <= "0000000000000000";
		mem(215)  <= "0000000000000000";
		mem(216)  <= "0000000000000000";
		mem(217)  <= "0000000000000000";
		mem(218)  <= "0000000000000000";
		mem(219)  <= "0000000000000000";
		mem(220)  <= "0000000000000000";
		mem(221)  <= "0000000000000000";
		mem(222)  <= "0000000000000000";
		mem(223)  <= "0000000000000000";
		mem(224)  <= "0000000000000000";
		mem(225)  <= "0000000000000000";
		mem(226)  <= "0000000000000000";
		mem(227)  <= "0000000000000000";
		mem(228)  <= "0000000000000000";
		mem(229)  <= "0000000000000000";
		mem(230)  <= "0000000000000000";
		mem(231)  <= "0000000000000000";
		mem(232)  <= "0000000000000000";
		mem(233)  <= "0000000000000000";
		mem(234)  <= "0000000000000000";
		mem(235)  <= "0000000000000000";
		mem(236)  <= "0000000000000000";
		mem(237)  <= "0000000000000000";
		mem(238)  <= "0000000000000000";
		mem(239)  <= "0000000000000000";
		mem(240)  <= "0000000000000000";
		mem(241)  <= "0000000000000000";
		mem(242)  <= "0000000000000000";
		mem(243)  <= "0000000000000000";
		mem(244)  <= "0000000000000000";
		mem(245)  <= "0000000000000000";
		mem(246)  <= "0000000000000000";
		mem(247)  <= "0000000000000000";
		mem(248)  <= "0000000000000000";
		mem(249)  <= "0000000000000000";
		mem(250)  <= "0000000000000000";
		mem(251)  <= "0000000000000000";
		mem(252)  <= "0000000000000000";
		mem(253)  <= "0000000000000000";
		mem(254)  <= "0000000000000000";
		mem(255)  <= "0000000000000000";
	else
	    -- read from memory
		if((leitura = '1'))then 
			saida_memoria(15 downto 0) <= mem(to_integer(unsigned(endereco_memoria)));
	-- write in memory		
		elsif ((escrita = '1')) then 		
			mem(to_integer(unsigned(endereco_memoria))) <= entrada_memoria(15 downto 0);
		end if;
	end if;		

						
end process;

end rtl;